--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   19:35:08 05/04/2019
-- Design Name:   
-- Module Name:   /home/aman/Desktop/IITB/CS226/project_ospf/CS226_OSPF/OSPF/lsup_tb2.vhd
-- Project Name:  OSPF
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: LSU_Parser
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY lsup_tb2 IS
END lsup_tb2;
 
ARCHITECTURE behavior OF lsup_tb2 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT LSU_Parser
    PORT(
         state_in : IN  std_logic_vector(3 downto 0);
         data_in : IN  std_logic_vector(7 downto 0);
         data_valid : IN  std_logic;
         clk : IN  std_logic;
         write_to_q : OUT  std_logic;
         qout : OUT  std_logic_vector(7 downto 0);
         ack_q_out : OUT  std_logic_vector(7 downto 0);
         ack_q_val : OUT  std_logic
        );
    END COMPONENT;
    COMPONENT Parser
    PORT(
         in1 : IN  std_logic_vector(7 downto 0);
         validity : IN  std_logic;
         clk : IN  std_logic;
         out1 : OUT  std_logic_vector(7 downto 0);
         hello_out : OUT  std_logic;
         ls_out : OUT  std_logic;
         telling_lsu : OUT  std_logic;
         telling_dd : OUT  std_logic;
         telling_plen : OUT  std_logic;
         telling_rid : OUT  std_logic;
         telling_lsr : OUT  std_logic;
         telling_neighbour : OUT  std_logic
        );
    END COMPONENT;

   --Inputs
   signal state_in : std_logic_vector(3 downto 0) := "0110";
   signal data_in : std_logic_vector(7 downto 0) := (others => '0');
   signal data_valid : std_logic := '0';
   signal clk : std_logic := '0';

 	--Outputs
   signal write_to_q : std_logic;
   signal qout : std_logic_vector(7 downto 0);
   signal ack_q_out : std_logic_vector(7 downto 0);
   signal ack_q_val : std_logic;
	signal in1 : std_logic_vector(7 downto 0);
	signal validity : std_logic;
	signal hello_out,ls_out : std_logic;
	signal telling : std_logic_vector(4 downto 0);
   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: LSU_Parser PORT MAP (
          state_in => state_in,
          data_in => data_in,
          data_valid => data_valid,
          clk => clk,
          write_to_q => write_to_q,
          qout => qout,
          ack_q_out => ack_q_out,
          ack_q_val => ack_q_val
        );
	uut1 : Parser PORT MAP (
			in1 => in1,
         validity => validity,
         clk => clk,
         out1 => data_in,
         hello_out => hello_out,
         ls_out => ls_out,
         telling_lsu => data_valid,
         telling_dd => telling(4),
         telling_plen => telling(3),
         telling_rid => telling(2),
         telling_lsr => telling(1),
         telling_neighbour => telling(0)
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		validity <= '1';
		in1 <= "00000000";
validity <= '1';
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00100000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "11011100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;



		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "01011100";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "11011100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000110";
		wait for clk_period;
		in1 <= "11001111";
		wait for clk_period;
		in1 <= "01100100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "01001000";
		wait for clk_period;
		in1 <= "11110011";
		wait for clk_period;
		in1 <= "11111100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00111100";
		wait for clk_period;
		in1 <= "10010011";
		wait for clk_period;
		in1 <= "00101111";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "01001000";
		wait for clk_period;

		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00100100";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;



		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "11101000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "01100100";
		wait for clk_period;
		in1 <= "10100101";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "01001000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00010100";
		wait for clk_period;
		in1 <= "00010100";
		wait for clk_period;
		in1 <= "00010100";
		wait for clk_period;
		in1 <= "00010100";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000111";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "10100110";
		wait for clk_period;
		in1 <= "01010000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00111100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00010101";
		wait for clk_period;
		in1 <= "11110000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000101";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "01001000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000010";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000100";
		wait for clk_period;
		in1 <= "00110010";
		wait for clk_period;
		in1 <= "00110010";
		wait for clk_period;
		in1 <= "00110010";
		wait for clk_period;
		in1 <= "00110010";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "11111111";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00001001";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000001";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000000";
		wait for clk_period;
		in1 <= "00000011";
		wait for clk_period;
		validity <= '0';
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
