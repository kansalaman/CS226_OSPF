LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
 
ENTITY tb_Main_Machine IS
END tb_Main_Machine;
 
ARCHITECTURE behavior OF tb_Main_Machine IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MainModule
    PORT(
         clk : IN  std_logic;
         in1 : IN  std_logic_vector(7 downto 0);
         in2 : IN  std_logic_vector(7 downto 0);
         in3 : IN  std_logic_vector(7 downto 0);
         in4 : IN  std_logic_vector(7 downto 0);
         in5 : IN  std_logic_vector(7 downto 0);
         in6 : IN  std_logic_vector(7 downto 0);
         in7 : IN  std_logic_vector(7 downto 0);
         in8 : IN  std_logic_vector(7 downto 0);
         in_val1 : IN  std_logic;
         in_val2 : IN  std_logic;
         in_val3 : IN  std_logic;
         in_val4 : IN  std_logic;
         in_val5 : IN  std_logic;
         in_val6 : IN  std_logic;
         in_val7 : IN  std_logic;
         in_val8 : IN  std_logic;
         out1 : OUT  std_logic_vector(7 downto 0);
         out2 : OUT  std_logic_vector(7 downto 0);
         out3 : OUT  std_logic_vector(7 downto 0);
         out4 : OUT  std_logic_vector(7 downto 0);
         out5 : OUT  std_logic_vector(7 downto 0);
         out6 : OUT  std_logic_vector(7 downto 0);
         out7 : OUT  std_logic_vector(7 downto 0);
         out8 : OUT  std_logic_vector(7 downto 0);
         out_val1 : OUT  std_logic;
         out_val2 : OUT std_logic;
         out_val3 : OUT std_logic;
         out_val4 : OUT std_logic;
         out_val5 : OUT std_logic;
         out_val6 : OUT std_logic;
         out_val7 : OUT std_logic;
         out_val8 : OUT std_logic
--         dijkstra_on : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal in1 : std_logic_vector(7 downto 0) := (others => '0');
   signal in2 : std_logic_vector(7 downto 0) := (others => '0');
   signal in3 : std_logic_vector(7 downto 0) := (others => '0');
   signal in4 : std_logic_vector(7 downto 0) := (others => '0');
   signal in5 : std_logic_vector(7 downto 0) := (others => '0');
   signal in6 : std_logic_vector(7 downto 0) := (others => '0');
   signal in7 : std_logic_vector(7 downto 0) := (others => '0');
   signal in8 : std_logic_vector(7 downto 0) := (others => '0');
   signal in_val1, in_val2, in_val3, in_val4, in_val5, in_val6, in_val7, in_val8 : std_logic:='0';
--   signal in_val2 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val3 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val4 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val5 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val6 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val7 : std_logic_vector(7 downto 0) := (others => '0');
--   signal in_val8 : std_logic_vector(7 downto 0) := (others => '0');
   signal out_val1 : std_logic := '0';
   signal out_val2 : std_logic := '0';
   signal out_val3 : std_logic := '0';
   signal out_val4 : std_logic := '0';
   signal out_val5 : std_logic := '0';
   signal out_val6 : std_logic := '0';
   signal out_val7 : std_logic := '0';
   signal out_val8 : std_logic := '0';
--   signal dijkstra_on : std_logic := '0';

 	--Outputs
   signal out1 : std_logic_vector(7 downto 0);
   signal out2 : std_logic_vector(7 downto 0);
   signal out3 : std_logic_vector(7 downto 0);
   signal out4 : std_logic_vector(7 downto 0);
   signal out5 : std_logic_vector(7 downto 0);
   signal out6 : std_logic_vector(7 downto 0);
   signal out7 : std_logic_vector(7 downto 0);
   signal out8 : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MainModule PORT MAP (
          clk => clk,
          in1 => in1,
          in2 => in2,
          in3 => in3,
          in4 => in4,
          in5 => in5,
          in6 => in6,
          in7 => in7,
          in8 => in8,
          in_val1 => in_val1,
          in_val2 => in_val2,
          in_val3 => in_val3,
          in_val4 => in_val4,
          in_val5 => in_val5,
          in_val6 => in_val6,
          in_val7 => in_val7,
          in_val8 => in_val8,
          out1 => out1,
          out2 => out2,
          out3 => out3,
          out4 => out4,
          out5 => out5,
          out6 => out6,
          out7 => out7,
          out8 => out8,
          out_val1 => out_val1,
          out_val2 => out_val2,
          out_val3 => out_val3,
          out_val4 => out_val4,
          out_val5 => out_val5,
          out_val6 => out_val6,
          out_val7 => out_val7,
          out_val8 => out_val8
--          dijkstra_on => dijkstra_on
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 95 ns;	
		
-- Sending Hello Packet from B at 95ns, using input port2
in_val2 <= '1';		
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00111000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="11101000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000111";
wait for clk_period;
in2<="11010000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
in_val2 <= '0';
wait for clk_period;

-- Sending Hello from C on port 3 after 50 cycles
wait for clk_period*50;

in_val3 <= '1';
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00111000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="11101000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000111";
wait for clk_period;
in3<="11010000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000000";
in_val3 <= '0';

-- Sending Empty DBD from B after 20 clk cycles
wait for clk_period*20;

in_val2 <= '1';
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00100000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="11011100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000111";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in_val2 <= '0';

-- Sending EMPTY DBD from C after 20 clock cycles

wait for 20*clk_period;

in_val3 <= '1';
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00100000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="11011100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000111";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00001010";
wait for clk_period;

in_val3 <= '0';

-- Reply DD_B after 200 clk_period 
wait for 200*clk_period;

in_val2 <= '1';
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="01011100";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="11011100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000110";
wait for clk_period;
in2<="00101000";
wait for clk_period;
in2<="01001010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="01001000";
wait for clk_period;
in2<="00110000";
wait for clk_period;
in2<="10010001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00111100";
wait for clk_period;
in2<="11010010";
wait for clk_period;
in2<="10010100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="01001000";
wait for clk_period;
in_val2 <= '0';

wait for 200*clk_period;
-- REPLY DBD FROM C after 200 clk cycles
in_val3 <= '1';
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="01011100";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="11011100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00001011";
wait for clk_period;
in3<="01001001";
wait for clk_period;
in3<="01111011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="01001000";
wait for clk_period;
in3<="11011100";
wait for clk_period;
in3<="00101011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00111100";
wait for clk_period;
in3<="10010100";
wait for clk_period;
in3<="00010000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="01001000";
wait for clk_period;
in_val3 <= '0';


-- LSR FROM B

wait for 120*clk_period;

in_val2 <= '1';
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00100100";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;

in_val2 <= '0';

-- SENDING LSR from C

wait for 300*clk_period;

in_val3 <= '1';
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00100100";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;

in_val3 <= '0';


-- Receiving LSU from B
wait for 50*clk_period;

in_val2 <= '1';
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2 <= "00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="11100101";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="11011111";
wait for clk_period;
in2<="01001111";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="01001000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00010100";
wait for clk_period;
in2<="00010100";
wait for clk_period;
in2<="00010100";
wait for clk_period;
in2<="00010100";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000111";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="10101010";
wait for clk_period;
in2<="11101110";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00111100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="10011010";
wait for clk_period;
in2<="00100111";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000101";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="01001000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000010";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000100";
wait for clk_period;
in2<="00110010";
wait for clk_period;
in2<="00110010";
wait for clk_period;
in2<="00110010";
wait for clk_period;
in2<="00110010";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="11111111";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00001001";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000011";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000001";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000000";
wait for clk_period;
in2<="00000011";
wait for clk_period;

in_val2 <= '0';


wait for 400*clk_period;

-- SENDING LSU from C
in_val3 <= '1';
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3 <= "00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="11100101";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="11010011";
wait for clk_period;
in3<="01011000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="01001000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00011110";
wait for clk_period;
in3<="00011110";
wait for clk_period;
in3<="00011110";
wait for clk_period;
in3<="00011110";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00001000";
wait for clk_period;
in3<="11011101";
wait for clk_period;
in3<="10001001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00111100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="01101010";
wait for clk_period;
in3<="00111110";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000101";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="01001000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000010";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000100";
wait for clk_period;
in3<="00110010";
wait for clk_period;
in3<="00110010";
wait for clk_period;
in3<="00110010";
wait for clk_period;
in3<="00110010";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="11111111";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00001001";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000011";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000001";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000000";
wait for clk_period;
in3<="00000011";
wait for clk_period;

in_val3 <= '0';


      wait;
   end process;

END;